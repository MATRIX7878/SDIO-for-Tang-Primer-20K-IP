LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SDDET IS
    PORT(DET : IN STD_LOGIC;
         LED : OUT STD_LOGIC
        );
END ENTITY;

ARCHITECTURE behavior OF SDDET IS

BEGIN
    PROCESS
        BEGIN
            WHILE DET LOOP
            END LOOP;
            LED <= '0';
    END PROCESS;
END ARCHITECTURE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SDCTRL IS

END ENTITY;

ARCHITECTURE Behavior OF SDCTRL IS
    COMPONENT SDDET IS
        PORT(DET : IN STD_LOGIC;
             LED : OUT STD_LOGIC
            );
    END COMPONENT;

    SIGNAL card : STD_LOGIC;

    BEGIN
        det : SDDET PORT MAP(DET => card);
   
END ARCHITECTURE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SDRW IS

END ENTITY;

ARCHITECTURE BEHAVIOR OF SDRW IS
    COMPONENT SDDET IS
        PORT(DET : IN STD_LOGIC;
             LED : OUT STD_LOGIC
            );
    END COMPONENT;

    SIGNAL card : STD_LOGIC;

    BEGIN
        det : SDDET PORT MAP(DET => card);
END ARCHITECTURE;