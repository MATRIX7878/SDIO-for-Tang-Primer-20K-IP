PACKAGE instructions IS
    TYPE SDCMDS IS (CMD0);
END PACKAGE;
