PACKAGE SDIOStates IS
    TYPE state IS (LOADDATA, SENDCMD, SENDDATA, READRESP, READDATA, DONE);
END PACKAGE;
